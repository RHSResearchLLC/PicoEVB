`include "sample_tests.vh"
